class AXI5_coverage extends uvm_component;

//=====================factory registration ============================

	`uvm_component_utils(AXI5_coverage)

//============================construction========================

	function new(string name="",uvm_component parent);
		super.new(name,parent);
	endfunction



endclass
